module decoder5_32(
    input [4:0] in,
    output [31:0] out
);

reg [31:0] out_reg;

always @(*) begin
    case (in)
        5'd0: out_reg = 32'b00000000000000000000000000000001;
        5'd1: out_reg = 32'b00000000000000000000000000000010;
        5'd2: out_reg = 32'b00000000000000000000000000000100;
        5'd3: out_reg = 32'b00000000000000000000000000001000;
        5'd4: out_reg = 32'b00000000000000000000000000010000;
        5'd5: out_reg = 32'b00000000000000000000000000100000;
        5'd6: out_reg = 32'b00000000000000000000000001000000;
        5'd7: out_reg = 32'b00000000000000000000000010000000;
        5'd8: out_reg = 32'b00000000000000000000000100000000;
        5'd9: out_reg = 32'b00000000000000000000001000000000;
        5'd10: out_reg = 32'b00000000000000000000010000000000;
        5'd11: out_reg = 32'b00000000000000000000100000000000;
        5'd12: out_reg = 32'b00000000000000000001000000000000;
        5'd13: out_reg = 32'b00000000000000000010000000000000;
        5'd14: out_reg = 32'b00000000000000000100000000000000;
        5'd15: out_reg = 32'b00000000000000001000000000000000;
        5'd16: out_reg = 32'b00000000000000010000000000000000;
        5'd17: out_reg = 32'b00000000000000100000000000000000;
        5'd18: out_reg = 32'b00000000000001000000000000000000;
        5'd19: out_reg = 32'b00000000000010000000000000000000;
        5'd20: out_reg = 32'b00000000000100000000000000000000;
        5'd21: out_reg = 32'b00000000001000000000000000000000;
        5'd22: out_reg = 32'b00000000010000000000000000000000;
        5'd23: out_reg = 32'b00000000100000000000000000000000;
        5'd24: out_reg = 32'b00000001000000000000000000000000;
        5'd25: out_reg = 32'b00000010000000000000000000000000;
        5'd26: out_reg = 32'b00000100000000000000000000000000;
        5'd27: out_reg = 32'b00001000000000000000000000000000;
        5'd28: out_reg = 32'b00010000000000000000000000000000;
        5'd29: out_reg = 32'b00100000000000000000000000000000;
        5'd30: out_reg = 32'b01000000000000000000000000000000;
        5'd31: out_reg = 32'b10000000000000000000000000000000;
        default: out_reg = 32'b00000000000000000000000000000000;
    endcase
end

assign out = out_reg;

endmodule